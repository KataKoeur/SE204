module reset (
  // port d'entrée
  input CLK,
  input NRST_in,
  // port de sortie
  output logic NRST_out
  );

parameter logic ACTIF_H = 1,



endmodule // reset
