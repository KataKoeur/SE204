module wshb_intercon (
  // interface
  wshb_if.slave  wshb_if_mire
  wshb_if.slave  wshb_if_vga
  wshb_if.master wshb_if_0
  );

endmodule // wshb_intercon
