module MED #(parameter SIZE = 8, NB_PIXEL = 9)(
        input [SIZE-1:0]DI,
        input logic DSI,
        input logic BYP,
        input logic CLK,
        output [SIZE-1:0]DO
        );



endmodule

