module foo();

initial
begin
	// $display est une tache système
	$display("hello world");
end

endmodule
