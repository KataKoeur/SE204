module MED #(parameter SIZE = 8)(
        input logic [SIZE-1:0]DI,
        input logic DSI,
        input logic nRST,
        input logic CLK,
        output logic [SIZE-1:0]DO,
        output logic DSO
        );


endmodule
