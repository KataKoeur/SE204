module mire (
  // mire interface
  wshb_if.master wshb_if_mire
  );

endmodule // mire
